library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.tfg_irene_package.ALL;
use IEEE.NUMERIC_STD.ALL;

entity VOT_INTERFAZ_ET2 is
Port ( 
		 dato_out_1 : in std_logic;
		 cero_1 : in std_logic;
		 dato_cero_1 : in std_logic;
		 padding_col2_1 : in std_logic;
		 padding_row2_1 : in std_logic;
		 col2_1 : in unsigned(log2c(column_size2 + 2*(conv2_padding)) - 1 downto 0);
		 p_row2_1: in unsigned( log2c(conv2_padding) downto 0); 
		 p_col2_1 : in unsigned( log2c(conv2_padding) downto 0);  
		 conv2_col_1 : in unsigned(log2c(conv2_column) - 1 downto 0);
		 conv2_fila_1 : in  unsigned(log2c(conv2_row) - 1 downto 0);
		 pool3_col_1 : in unsigned(log2c(pool3_column) - 1 downto 0);
		 pool3_fila_1 : in  unsigned(log2c(pool3_row) - 1 downto 0);
		 dato_out_2 : in std_logic;
		 cero_2 : in std_logic;
		 dato_cero_2 : in std_logic;
		 padding_col2_2 : in std_logic;
		 padding_row2_2 : in std_logic;
		 col2_2 : in unsigned(log2c(column_size2 + 2*(conv2_padding)) - 1 downto 0);
		 p_row2_2: in unsigned( log2c(conv2_padding) downto 0); 
		 p_col2_2 : in unsigned( log2c(conv2_padding) downto 0);  
		 conv2_col_2 : in unsigned(log2c(conv2_column) - 1 downto 0);
		 conv2_fila_2 : in  unsigned(log2c(conv2_row) - 1 downto 0);
		 pool3_col_2 : in unsigned(log2c(pool3_column) - 1 downto 0);
		 pool3_fila_2 : in  unsigned(log2c(pool3_row) - 1 downto 0);
		 dato_out_3 : in std_logic;
		 cero_3 : in std_logic;
		 dato_cero_3 : in std_logic;
		 padding_col2_3 : in std_logic;
		 padding_row2_3 : in std_logic;
		 col2_3 : in unsigned(log2c(column_size2 + 2*(conv2_padding)) - 1 downto 0);
		 p_row2_3: in unsigned( log2c(conv2_padding) downto 0); 
		 p_col2_3 : in unsigned( log2c(conv2_padding) downto 0);  
		 conv2_col_3 : in unsigned(log2c(conv2_column) - 1 downto 0);
		 conv2_fila_3 : in  unsigned(log2c(conv2_row) - 1 downto 0);
		 pool3_col_3 : in unsigned(log2c(pool3_column) - 1 downto 0);
		 pool3_fila_3 : in  unsigned(log2c(pool3_row) - 1 downto 0);
		 dato_out_v : out std_logic;
		 cero_v : out std_logic;
		 dato_cero_v : out std_logic;
		 padding_col2_v : out std_logic;
		 padding_row2_v : out std_logic;
		 col2_v : out unsigned(log2c(column_size2 + 2*(conv2_padding)) - 1 downto 0);
		 p_row2_v: out unsigned( log2c(conv2_padding) downto 0); 
		 p_col2_v : out unsigned( log2c(conv2_padding) downto 0);  
		 conv2_col_v : out unsigned(log2c(conv2_column) - 1 downto 0);
		 conv2_fila_v : out  unsigned(log2c(conv2_row) - 1 downto 0);
		 pool3_col_v : out unsigned(log2c(pool3_column) - 1 downto 0);
		 pool3_fila_v : out  unsigned(log2c(pool3_row) - 1 downto 0));
end VOT_Interfaz_ET2;
architecture Behavioral of VOT_Interfaz_ET2 is
begin
dato_out_v <= (dato_out_1 and dato_out_2) or (dato_out_1 and dato_out_3) or (dato_out_2 and dato_out_3);
cero_v <= (cero_1 and cero_2) or (cero_1 and cero_3) or (cero_2 and cero_3);
dato_cero_v <= (dato_cero_1 and dato_cero_2) or (dato_cero_1 and dato_cero_3) or (dato_cero_2 and dato_cero_3);
		 padding_col2_v <= (padding_col2_1 and padding_col2_2) or (padding_col2_1 and padding_col2_3) or (padding_col2_2 and padding_col2_3);
		 padding_row2_v <= (padding_row2_1 and padding_row2_2) or (padding_row2_1 and padding_row2_3) or (padding_row2_2 and padding_row2_3);
		 col2_v <= (col2_1 and col2_2) or (col2_1 and col2_3) or (col2_2 and col2_3);
		 p_row2_v <= (p_row2_1 and p_row2_2) or (p_row2_1 and p_row2_3) or (p_row2_2 and p_row2_3);
		 p_col2_v <= (p_col2_1 and p_col2_2) or (p_col2_1 and p_col2_3) or (p_col2_2 and p_col2_3);  
		 conv2_col_v <= (conv2_col_1 and conv2_col_2) or (conv2_col_1 and conv2_col_3) or (conv2_col_2 and conv2_col_3);
		 conv2_fila_v <= (conv2_fila_1 and conv2_fila_2) or (conv2_fila_1 and conv2_fila_3) or (conv2_fila_2 and conv2_fila_3);
		 pool3_col_v <= (pool3_col_1 and pool3_col_2) or (pool3_col_1 and pool3_col_3) or (pool3_col_2 and pool3_col_3);
		 pool3_fila_v <= (pool3_fila_1 and pool3_fila_2) or (pool3_fila_1 and pool3_fila_3) or (pool3_fila_2 and pool3_fila_3);
end Behavioral;
