library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.tfg_irene_package.ALL;
use IEEE.NUMERIC_STD.ALL;

entity VOT_Register_FCL2 is
    Port (  
       data_out_1 : in vector_L2fc_activations(0 to number_of_inputs_L3fc-1);
       data_out_2 : in vector_L2fc_activations(0 to number_of_inputs_L3fc-1);
       data_out_3 : in vector_L2fc_activations(0 to number_of_inputs_L3fc-1);
       data_out_v : out vector_L2fc_activations(0 to number_of_inputs_L3fc-1));
end VOT_Register_FCL2;

architecture Behavioral of VOT_Register_FCL2 is

begin

data_out_v(0) <= (data_out_1(0) and data_out_2(0)) or (data_out_1(0) and data_out_3(0)) or (data_out_2(0) and data_out_3(0));
data_out_v(1) <= (data_out_1(1) and data_out_2(1)) or (data_out_1(1) and data_out_3(1)) or (data_out_2(1) and data_out_3(1));
data_out_v(2) <= (data_out_1(2) and data_out_2(2)) or (data_out_1(2) and data_out_3(2)) or (data_out_2(2) and data_out_3(2));
data_out_v(3) <= (data_out_1(3) and data_out_2(3)) or (data_out_1(3) and data_out_3(3)) or (data_out_2(3) and data_out_3(3));
data_out_v(4) <= (data_out_1(4) and data_out_2(4)) or (data_out_1(4) and data_out_3(4)) or (data_out_2(4) and data_out_3(4));
data_out_v(5) <= (data_out_1(5) and data_out_2(5)) or (data_out_1(5) and data_out_3(5)) or (data_out_2(5) and data_out_3(5));
data_out_v(6) <= (data_out_1(6) and data_out_2(6)) or (data_out_1(6) and data_out_3(6)) or (data_out_2(6) and data_out_3(6));
data_out_v(7) <= (data_out_1(7) and data_out_2(7)) or (data_out_1(7) and data_out_3(7)) or (data_out_2(7) and data_out_3(7));
data_out_v(8) <= (data_out_1(8) and data_out_2(8)) or (data_out_1(8) and data_out_3(8)) or (data_out_2(8) and data_out_3(8));
data_out_v(9) <= (data_out_1(9) and data_out_2(9)) or (data_out_1(9) and data_out_3(9)) or (data_out_2(9) and data_out_3(9));
data_out_v(10) <= (data_out_1(10) and data_out_2(10)) or (data_out_1(10) and data_out_3(10)) or (data_out_2(10) and data_out_3(10));
data_out_v(11) <= (data_out_1(11) and data_out_2(11)) or (data_out_1(11) and data_out_3(11)) or (data_out_2(11) and data_out_3(11));
data_out_v(12) <= (data_out_1(12) and data_out_2(12)) or (data_out_1(12) and data_out_3(12)) or (data_out_2(12) and data_out_3(12));
data_out_v(13) <= (data_out_1(13) and data_out_2(13)) or (data_out_1(13) and data_out_3(13)) or (data_out_2(13) and data_out_3(13));
data_out_v(14) <= (data_out_1(14) and data_out_2(14)) or (data_out_1(14) and data_out_3(14)) or (data_out_2(14) and data_out_3(14));
data_out_v(15) <= (data_out_1(15) and data_out_2(15)) or (data_out_1(15) and data_out_3(15)) or (data_out_2(15) and data_out_3(15));
data_out_v(16) <= (data_out_1(16) and data_out_2(16)) or (data_out_1(16) and data_out_3(16)) or (data_out_2(16) and data_out_3(16));
data_out_v(17) <= (data_out_1(17) and data_out_2(17)) or (data_out_1(17) and data_out_3(17)) or (data_out_2(17) and data_out_3(17));
data_out_v(18) <= (data_out_1(18) and data_out_2(18)) or (data_out_1(18) and data_out_3(18)) or (data_out_2(18) and data_out_3(18));
data_out_v(19) <= (data_out_1(19) and data_out_2(19)) or (data_out_1(19) and data_out_3(19)) or (data_out_2(19) and data_out_3(19));
data_out_v(20) <= (data_out_1(20) and data_out_2(20)) or (data_out_1(20) and data_out_3(20)) or (data_out_2(20) and data_out_3(20));
data_out_v(21) <= (data_out_1(21) and data_out_2(21)) or (data_out_1(21) and data_out_3(21)) or (data_out_2(21) and data_out_3(21));
data_out_v(22) <= (data_out_1(22) and data_out_2(22)) or (data_out_1(22) and data_out_3(22)) or (data_out_2(22) and data_out_3(22));
data_out_v(23) <= (data_out_1(23) and data_out_2(23)) or (data_out_1(23) and data_out_3(23)) or (data_out_2(23) and data_out_3(23));
data_out_v(24) <= (data_out_1(24) and data_out_2(24)) or (data_out_1(24) and data_out_3(24)) or (data_out_2(24) and data_out_3(24));
data_out_v(25) <= (data_out_1(25) and data_out_2(25)) or (data_out_1(25) and data_out_3(25)) or (data_out_2(25) and data_out_3(25));
data_out_v(26) <= (data_out_1(26) and data_out_2(26)) or (data_out_1(26) and data_out_3(26)) or (data_out_2(26) and data_out_3(26));
data_out_v(27) <= (data_out_1(27) and data_out_2(27)) or (data_out_1(27) and data_out_3(27)) or (data_out_2(27) and data_out_3(27));
data_out_v(28) <= (data_out_1(28) and data_out_2(28)) or (data_out_1(28) and data_out_3(28)) or (data_out_2(28) and data_out_3(28));
data_out_v(29) <= (data_out_1(29) and data_out_2(29)) or (data_out_1(29) and data_out_3(29)) or (data_out_2(29) and data_out_3(29));
data_out_v(30) <= (data_out_1(30) and data_out_2(30)) or (data_out_1(30) and data_out_3(30)) or (data_out_2(30) and data_out_3(30));
data_out_v(31) <= (data_out_1(31) and data_out_2(31)) or (data_out_1(31) and data_out_3(31)) or (data_out_2(31) and data_out_3(31));
data_out_v(32) <= (data_out_1(32) and data_out_2(32)) or (data_out_1(32) and data_out_3(32)) or (data_out_2(32) and data_out_3(32));
data_out_v(33) <= (data_out_1(33) and data_out_2(33)) or (data_out_1(33) and data_out_3(33)) or (data_out_2(33) and data_out_3(33));
data_out_v(34) <= (data_out_1(34) and data_out_2(34)) or (data_out_1(34) and data_out_3(34)) or (data_out_2(34) and data_out_3(34));
data_out_v(35) <= (data_out_1(35) and data_out_2(35)) or (data_out_1(35) and data_out_3(35)) or (data_out_2(35) and data_out_3(35));
data_out_v(36) <= (data_out_1(36) and data_out_2(36)) or (data_out_1(36) and data_out_3(36)) or (data_out_2(36) and data_out_3(36));
data_out_v(37) <= (data_out_1(37) and data_out_2(37)) or (data_out_1(37) and data_out_3(37)) or (data_out_2(37) and data_out_3(37));
data_out_v(38) <= (data_out_1(38) and data_out_2(38)) or (data_out_1(38) and data_out_3(38)) or (data_out_2(38) and data_out_3(38));
data_out_v(39) <= (data_out_1(39) and data_out_2(39)) or (data_out_1(39) and data_out_3(39)) or (data_out_2(39) and data_out_3(39));
data_out_v(40) <= (data_out_1(40) and data_out_2(40)) or (data_out_1(40) and data_out_3(40)) or (data_out_2(40) and data_out_3(40));
data_out_v(41) <= (data_out_1(41) and data_out_2(41)) or (data_out_1(41) and data_out_3(41)) or (data_out_2(41) and data_out_3(41));
data_out_v(42) <= (data_out_1(42) and data_out_2(42)) or (data_out_1(42) and data_out_3(42)) or (data_out_2(42) and data_out_3(42));
data_out_v(43) <= (data_out_1(43) and data_out_2(43)) or (data_out_1(43) and data_out_3(43)) or (data_out_2(43) and data_out_3(43));
data_out_v(44) <= (data_out_1(44) and data_out_2(44)) or (data_out_1(44) and data_out_3(44)) or (data_out_2(44) and data_out_3(44));
data_out_v(45) <= (data_out_1(45) and data_out_2(45)) or (data_out_1(45) and data_out_3(45)) or (data_out_2(45) and data_out_3(45));
data_out_v(46) <= (data_out_1(46) and data_out_2(46)) or (data_out_1(46) and data_out_3(46)) or (data_out_2(46) and data_out_3(46));
data_out_v(47) <= (data_out_1(47) and data_out_2(47)) or (data_out_1(47) and data_out_3(47)) or (data_out_2(47) and data_out_3(47));
data_out_v(48) <= (data_out_1(48) and data_out_2(48)) or (data_out_1(48) and data_out_3(48)) or (data_out_2(48) and data_out_3(48));
data_out_v(49) <= (data_out_1(49) and data_out_2(49)) or (data_out_1(49) and data_out_3(49)) or (data_out_2(49) and data_out_3(49));
data_out_v(50) <= (data_out_1(50) and data_out_2(50)) or (data_out_1(50) and data_out_3(50)) or (data_out_2(50) and data_out_3(50));
data_out_v(51) <= (data_out_1(51) and data_out_2(51)) or (data_out_1(51) and data_out_3(51)) or (data_out_2(51) and data_out_3(51));
data_out_v(52) <= (data_out_1(52) and data_out_2(52)) or (data_out_1(52) and data_out_3(52)) or (data_out_2(52) and data_out_3(52));
data_out_v(53) <= (data_out_1(53) and data_out_2(53)) or (data_out_1(53) and data_out_3(53)) or (data_out_2(53) and data_out_3(53));
data_out_v(54) <= (data_out_1(54) and data_out_2(54)) or (data_out_1(54) and data_out_3(54)) or (data_out_2(54) and data_out_3(54));
data_out_v(55) <= (data_out_1(55) and data_out_2(55)) or (data_out_1(55) and data_out_3(55)) or (data_out_2(55) and data_out_3(55));
data_out_v(56) <= (data_out_1(56) and data_out_2(56)) or (data_out_1(56) and data_out_3(56)) or (data_out_2(56) and data_out_3(56));
data_out_v(57) <= (data_out_1(57) and data_out_2(57)) or (data_out_1(57) and data_out_3(57)) or (data_out_2(57) and data_out_3(57));
data_out_v(58) <= (data_out_1(58) and data_out_2(58)) or (data_out_1(58) and data_out_3(58)) or (data_out_2(58) and data_out_3(58));
data_out_v(59) <= (data_out_1(59) and data_out_2(59)) or (data_out_1(59) and data_out_3(59)) or (data_out_2(59) and data_out_3(59));
data_out_v(60) <= (data_out_1(60) and data_out_2(60)) or (data_out_1(60) and data_out_3(60)) or (data_out_2(60) and data_out_3(60));
data_out_v(61) <= (data_out_1(61) and data_out_2(61)) or (data_out_1(61) and data_out_3(61)) or (data_out_2(61) and data_out_3(61));
data_out_v(62) <= (data_out_1(62) and data_out_2(62)) or (data_out_1(62) and data_out_3(62)) or (data_out_2(62) and data_out_3(62));
data_out_v(63) <= (data_out_1(63) and data_out_2(63)) or (data_out_1(63) and data_out_3(63)) or (data_out_2(63) and data_out_3(63));
data_out_v(64) <= (data_out_1(64) and data_out_2(64)) or (data_out_1(64) and data_out_3(64)) or (data_out_2(64) and data_out_3(64));
data_out_v(65) <= (data_out_1(65) and data_out_2(65)) or (data_out_1(65) and data_out_3(65)) or (data_out_2(65) and data_out_3(65));
data_out_v(66) <= (data_out_1(66) and data_out_2(66)) or (data_out_1(66) and data_out_3(66)) or (data_out_2(66) and data_out_3(66));
data_out_v(67) <= (data_out_1(67) and data_out_2(67)) or (data_out_1(67) and data_out_3(67)) or (data_out_2(67) and data_out_3(67));
data_out_v(68) <= (data_out_1(68) and data_out_2(68)) or (data_out_1(68) and data_out_3(68)) or (data_out_2(68) and data_out_3(68));
data_out_v(69) <= (data_out_1(69) and data_out_2(69)) or (data_out_1(69) and data_out_3(69)) or (data_out_2(69) and data_out_3(69));
data_out_v(70) <= (data_out_1(70) and data_out_2(70)) or (data_out_1(70) and data_out_3(70)) or (data_out_2(70) and data_out_3(70));
data_out_v(71) <= (data_out_1(71) and data_out_2(71)) or (data_out_1(71) and data_out_3(71)) or (data_out_2(71) and data_out_3(71));
data_out_v(72) <= (data_out_1(72) and data_out_2(72)) or (data_out_1(72) and data_out_3(72)) or (data_out_2(72) and data_out_3(72));
data_out_v(73) <= (data_out_1(73) and data_out_2(73)) or (data_out_1(73) and data_out_3(73)) or (data_out_2(73) and data_out_3(73));
data_out_v(74) <= (data_out_1(74) and data_out_2(74)) or (data_out_1(74) and data_out_3(74)) or (data_out_2(74) and data_out_3(74));
data_out_v(75) <= (data_out_1(75) and data_out_2(75)) or (data_out_1(75) and data_out_3(75)) or (data_out_2(75) and data_out_3(75));
data_out_v(76) <= (data_out_1(76) and data_out_2(76)) or (data_out_1(76) and data_out_3(76)) or (data_out_2(76) and data_out_3(76));
data_out_v(77) <= (data_out_1(77) and data_out_2(77)) or (data_out_1(77) and data_out_3(77)) or (data_out_2(77) and data_out_3(77));
data_out_v(78) <= (data_out_1(78) and data_out_2(78)) or (data_out_1(78) and data_out_3(78)) or (data_out_2(78) and data_out_3(78));
data_out_v(79) <= (data_out_1(79) and data_out_2(79)) or (data_out_1(79) and data_out_3(79)) or (data_out_2(79) and data_out_3(79));
data_out_v(80) <= (data_out_1(80) and data_out_2(80)) or (data_out_1(80) and data_out_3(80)) or (data_out_2(80) and data_out_3(80));
data_out_v(81) <= (data_out_1(81) and data_out_2(81)) or (data_out_1(81) and data_out_3(81)) or (data_out_2(81) and data_out_3(81));
data_out_v(82) <= (data_out_1(82) and data_out_2(82)) or (data_out_1(82) and data_out_3(82)) or (data_out_2(82) and data_out_3(82));
data_out_v(83) <= (data_out_1(83) and data_out_2(83)) or (data_out_1(83) and data_out_3(83)) or (data_out_2(83) and data_out_3(83));
end Behavioral;
