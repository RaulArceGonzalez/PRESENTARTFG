--Image5 is 5 predicted 5;
LIBRARY IEEE;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE work.tfg_irene_package.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.MATH_REAL.ALL;
ENTITY Mock_Memory IS
	PORT (
		clk : IN STD_LOGIC;
		rst : IN STD_LOGIC;
		address : IN STD_LOGIC_VECTOR(log2c(number_of_inputs) - 1 DOWNTO 0);
		data_out : OUT STD_LOGIC_VECTOR(input_sizeL1 - 1 DOWNTO 0));
END Mock_Memory;
ARCHITECTURE Behavioral OF Mock_Memory IS
	SIGNAL data_out_next, data_out_reg : STD_LOGIC_VECTOR(input_sizeL1 - 1 DOWNTO 0);
BEGIN
	PROCESS (clk)
	BEGIN
		IF rising_edge(clk) THEN
			IF (rst = '0') THEN
				data_out_reg <= (OTHERS => '0');
			ELSE
				data_out_reg <= data_out_next;
			END IF;
		END IF;
	END PROCESS;
	WITH address SELECT data_out_next <=
		"00000000" WHEN "0000000000", -- 0
		"00000000" WHEN "0000000001", -- 1
		"00000000" WHEN "0000000010", -- 2
		"00000000" WHEN "0000000011", -- 3
		"00000000" WHEN "0000000100", -- 4
		"00000000" WHEN "0000000101", -- 5
		"00000000" WHEN "0000000110", -- 6
		"00000000" WHEN "0000000111", -- 7
		"00000000" WHEN "0000001000", -- 8
		"00000000" WHEN "0000001001", -- 9
		"00000000" WHEN "0000001010", -- 10
		"00000000" WHEN "0000001011", -- 11
		"00000000" WHEN "0000001100", -- 12
		"00000000" WHEN "0000001101", -- 13
		"00000000" WHEN "0000001110", -- 14
		"00000000" WHEN "0000001111", -- 15
		"00000000" WHEN "0000010000", -- 16
		"00000000" WHEN "0000010001", -- 17
		"00000000" WHEN "0000010010", -- 18
		"00000000" WHEN "0000010011", -- 19
		"00000000" WHEN "0000010100", -- 20
		"00000000" WHEN "0000010101", -- 21
		"00000000" WHEN "0000010110", -- 22
		"00000000" WHEN "0000010111", -- 23
		"00000000" WHEN "0000011000", -- 24
		"00000000" WHEN "0000011001", -- 25
		"00000000" WHEN "0000011010", -- 26
		"00000000" WHEN "0000011011", -- 27
		"00000000" WHEN "0000011100", -- 28
		"00000000" WHEN "0000011101", -- 29
		"00000000" WHEN "0000011110", -- 30
		"00000000" WHEN "0000011111", -- 31
		"00000000" WHEN "0000100000", -- 32
		"00000000" WHEN "0000100001", -- 33
		"00000000" WHEN "0000100010", -- 34
		"00000000" WHEN "0000100011", -- 35
		"00000000" WHEN "0000100100", -- 36
		"00000000" WHEN "0000100101", -- 37
		"00000000" WHEN "0000100110", -- 38
		"00000000" WHEN "0000100111", -- 39
		"00000000" WHEN "0000101000", -- 40
		"00000000" WHEN "0000101001", -- 41
		"00000000" WHEN "0000101010", -- 42
		"00000000" WHEN "0000101011", -- 43
		"00000000" WHEN "0000101100", -- 44
		"00000000" WHEN "0000101101", -- 45
		"00000000" WHEN "0000101110", -- 46
		"00000000" WHEN "0000101111", -- 47
		"00000000" WHEN "0000110000", -- 48
		"00000000" WHEN "0000110001", -- 49
		"00000000" WHEN "0000110010", -- 50
		"00000000" WHEN "0000110011", -- 51
		"00000000" WHEN "0000110100", -- 52
		"00000000" WHEN "0000110101", -- 53
		"00000000" WHEN "0000110110", -- 54
		"00000000" WHEN "0000110111", -- 55
		"00000000" WHEN "0000111000", -- 56
		"00000000" WHEN "0000111001", -- 57
		"00000000" WHEN "0000111010", -- 58
		"00000000" WHEN "0000111011", -- 59
		"00000000" WHEN "0000111100", -- 60
		"00000000" WHEN "0000111101", -- 61
		"00000000" WHEN "0000111110", -- 62
		"00000000" WHEN "0000111111", -- 63
		"00000000" WHEN "0001000000", -- 64
		"00000000" WHEN "0001000001", -- 65
		"00000000" WHEN "0001000010", -- 66
		"00000000" WHEN "0001000011", -- 67
		"00000000" WHEN "0001000100", -- 68
		"00000000" WHEN "0001000101", -- 69
		"00000000" WHEN "0001000110", -- 70
		"00000000" WHEN "0001000111", -- 71
		"00000000" WHEN "0001001000", -- 72
		"00000000" WHEN "0001001001", -- 73
		"00000000" WHEN "0001001010", -- 74
		"00000000" WHEN "0001001011", -- 75
		"00000000" WHEN "0001001100", -- 76
		"00000000" WHEN "0001001101", -- 77
		"00000000" WHEN "0001001110", -- 78
		"00000000" WHEN "0001001111", -- 79
		"00000000" WHEN "0001010000", -- 80
		"00000000" WHEN "0001010001", -- 81
		"00000000" WHEN "0001010010", -- 82
		"00000000" WHEN "0001010011", -- 83
		"00000000" WHEN "0001010100", -- 84
		"00000000" WHEN "0001010101", -- 85
		"00000000" WHEN "0001010110", -- 86
		"00000000" WHEN "0001010111", -- 87
		"00000000" WHEN "0001011000", -- 88
		"00000000" WHEN "0001011001", -- 89
		"00000000" WHEN "0001011010", -- 90
		"00000000" WHEN "0001011011", -- 91
		"00000000" WHEN "0001011100", -- 92
		"00000000" WHEN "0001011101", -- 93
		"00000000" WHEN "0001011110", -- 94
		"00000000" WHEN "0001011111", -- 95
		"00000000" WHEN "0001100000", -- 96
		"00000000" WHEN "0001100001", -- 97
		"00000000" WHEN "0001100010", -- 98
		"00000000" WHEN "0001100011", -- 99
		"00000000" WHEN "0001100100", -- 100
		"00000000" WHEN "0001100101", -- 101
		"00000000" WHEN "0001100110", -- 102
		"00000000" WHEN "0001100111", -- 103
		"00000000" WHEN "0001101000", -- 104
		"00000000" WHEN "0001101001", -- 105
		"00000000" WHEN "0001101010", -- 106
		"00000000" WHEN "0001101011", -- 107
		"00000000" WHEN "0001101100", -- 108
		"00000000" WHEN "0001101101", -- 109
		"00000000" WHEN "0001101110", -- 110
		"00000000" WHEN "0001101111", -- 111
		"00000000" WHEN "0001110000", -- 112
		"00000000" WHEN "0001110001", -- 113
		"00000000" WHEN "0001110010", -- 114
		"00000000" WHEN "0001110011", -- 115
		"00000000" WHEN "0001110100", -- 116
		"00000000" WHEN "0001110101", -- 117
		"00000000" WHEN "0001110110", -- 118
		"00000000" WHEN "0001110111", -- 119
		"00000000" WHEN "0001111000", -- 120
		"00000000" WHEN "0001111001", -- 121
		"00000000" WHEN "0001111010", -- 122
		"00000000" WHEN "0001111011", -- 123
		"00000000" WHEN "0001111100", -- 124
		"00000000" WHEN "0001111101", -- 125
		"00000000" WHEN "0001111110", -- 126
		"00000000" WHEN "0001111111", -- 127
		"00000000" WHEN "0010000000", -- 128
		"00000000" WHEN "0010000001", -- 129
		"00000000" WHEN "0010000010", -- 130
		"00000000" WHEN "0010000011", -- 131
		"00000000" WHEN "0010000100", -- 132
		"00000000" WHEN "0010000101", -- 133
		"00000000" WHEN "0010000110", -- 134
		"00000000" WHEN "0010000111", -- 135
		"00000000" WHEN "0010001000", -- 136
		"00000000" WHEN "0010001001", -- 137
		"00000000" WHEN "0010001010", -- 138
		"00000000" WHEN "0010001011", -- 139
		"00000000" WHEN "0010001100", -- 140
		"00000000" WHEN "0010001101", -- 141
		"00000000" WHEN "0010001110", -- 142
		"00000000" WHEN "0010001111", -- 143
		"00000000" WHEN "0010010000", -- 144
		"00000000" WHEN "0010010001", -- 145
		"00000000" WHEN "0010010010", -- 146
		"00000000" WHEN "0010010011", -- 147
		"00000000" WHEN "0010010100", -- 148
		"00000000" WHEN "0010010101", -- 149
		"00000000" WHEN "0010010110", -- 150
		"00000000" WHEN "0010010111", -- 151
		"00000000" WHEN "0010011000", -- 152
		"00000100" WHEN "0010011001", -- 153
		"00000100" WHEN "0010011010", -- 154
		"00000100" WHEN "0010011011", -- 155
		"00011111" WHEN "0010011100", -- 156
		"00100010" WHEN "0010011101", -- 157
		"00101011" WHEN "0010011110", -- 158
		"00000110" WHEN "0010011111", -- 159
		"00101001" WHEN "0010100000", -- 160
		"01000000" WHEN "0010100001", -- 161
		"00111101" WHEN "0010100010", -- 162
		"00011111" WHEN "0010100011", -- 163
		"00000000" WHEN "0010100100", -- 164
		"00000000" WHEN "0010100101", -- 165
		"00000000" WHEN "0010100110", -- 166
		"00000000" WHEN "0010100111", -- 167
		"00000000" WHEN "0010101000", -- 168
		"00000000" WHEN "0010101001", -- 169
		"00000000" WHEN "0010101010", -- 170
		"00000000" WHEN "0010101011", -- 171
		"00000000" WHEN "0010101100", -- 172
		"00000000" WHEN "0010101101", -- 173
		"00000000" WHEN "0010101110", -- 174
		"00000000" WHEN "0010101111", -- 175
		"00000111" WHEN "0010110000", -- 176
		"00001001" WHEN "0010110001", -- 177
		"00010111" WHEN "0010110010", -- 178
		"00100110" WHEN "0010110011", -- 179
		"00101010" WHEN "0010110100", -- 180
		"00111111" WHEN "0010110101", -- 181
		"00111111" WHEN "0010110110", -- 182
		"00111111" WHEN "0010110111", -- 183
		"00111111" WHEN "0010111000", -- 184
		"00111111" WHEN "0010111001", -- 185
		"00111000" WHEN "0010111010", -- 186
		"00101011" WHEN "0010111011", -- 187
		"00111111" WHEN "0010111100", -- 188
		"00111100" WHEN "0010111101", -- 189
		"00110000" WHEN "0010111110", -- 190
		"00010000" WHEN "0010111111", -- 191
		"00000000" WHEN "0011000000", -- 192
		"00000000" WHEN "0011000001", -- 193
		"00000000" WHEN "0011000010", -- 194
		"00000000" WHEN "0011000011", -- 195
		"00000000" WHEN "0011000100", -- 196
		"00000000" WHEN "0011000101", -- 197
		"00000000" WHEN "0011000110", -- 198
		"00000000" WHEN "0011000111", -- 199
		"00000000" WHEN "0011001000", -- 200
		"00000000" WHEN "0011001001", -- 201
		"00000000" WHEN "0011001010", -- 202
		"00001100" WHEN "0011001011", -- 203
		"00111011" WHEN "0011001100", -- 204
		"00111111" WHEN "0011001101", -- 205
		"00111111" WHEN "0011001110", -- 206
		"00111111" WHEN "0011001111", -- 207
		"00111111" WHEN "0011010000", -- 208
		"00111111" WHEN "0011010001", -- 209
		"00111111" WHEN "0011010010", -- 210
		"00111111" WHEN "0011010011", -- 211
		"00111111" WHEN "0011010100", -- 212
		"00111110" WHEN "0011010101", -- 213
		"00010111" WHEN "0011010110", -- 214
		"00010100" WHEN "0011010111", -- 215
		"00010100" WHEN "0011011000", -- 216
		"00001110" WHEN "0011011001", -- 217
		"00001001" WHEN "0011011010", -- 218
		"00000000" WHEN "0011011011", -- 219
		"00000000" WHEN "0011011100", -- 220
		"00000000" WHEN "0011011101", -- 221
		"00000000" WHEN "0011011110", -- 222
		"00000000" WHEN "0011011111", -- 223
		"00000000" WHEN "0011100000", -- 224
		"00000000" WHEN "0011100001", -- 225
		"00000000" WHEN "0011100010", -- 226
		"00000000" WHEN "0011100011", -- 227
		"00000000" WHEN "0011100100", -- 228
		"00000000" WHEN "0011100101", -- 229
		"00000000" WHEN "0011100110", -- 230
		"00000100" WHEN "0011100111", -- 231
		"00110110" WHEN "0011101000", -- 232
		"00111111" WHEN "0011101001", -- 233
		"00111111" WHEN "0011101010", -- 234
		"00111111" WHEN "0011101011", -- 235
		"00111111" WHEN "0011101100", -- 236
		"00111111" WHEN "0011101101", -- 237
		"00110001" WHEN "0011101110", -- 238
		"00101101" WHEN "0011101111", -- 239
		"00111101" WHEN "0011110000", -- 240
		"00111100" WHEN "0011110001", -- 241
		"00000000" WHEN "0011110010", -- 242
		"00000000" WHEN "0011110011", -- 243
		"00000000" WHEN "0011110100", -- 244
		"00000000" WHEN "0011110101", -- 245
		"00000000" WHEN "0011110110", -- 246
		"00000000" WHEN "0011110111", -- 247
		"00000000" WHEN "0011111000", -- 248
		"00000000" WHEN "0011111001", -- 249
		"00000000" WHEN "0011111010", -- 250
		"00000000" WHEN "0011111011", -- 251
		"00000000" WHEN "0011111100", -- 252
		"00000000" WHEN "0011111101", -- 253
		"00000000" WHEN "0011111110", -- 254
		"00000000" WHEN "0011111111", -- 255
		"00000000" WHEN "0100000000", -- 256
		"00000000" WHEN "0100000001", -- 257
		"00000000" WHEN "0100000010", -- 258
		"00000000" WHEN "0100000011", -- 259
		"00010100" WHEN "0100000100", -- 260
		"00100111" WHEN "0100000101", -- 261
		"00011010" WHEN "0100000110", -- 262
		"00111111" WHEN "0100000111", -- 263
		"00111111" WHEN "0100001000", -- 264
		"00110011" WHEN "0100001001", -- 265
		"00000010" WHEN "0100001010", -- 266
		"00000000" WHEN "0100001011", -- 267
		"00001010" WHEN "0100001100", -- 268
		"00100110" WHEN "0100001101", -- 269
		"00000000" WHEN "0100001110", -- 270
		"00000000" WHEN "0100001111", -- 271
		"00000000" WHEN "0100010000", -- 272
		"00000000" WHEN "0100010001", -- 273
		"00000000" WHEN "0100010010", -- 274
		"00000000" WHEN "0100010011", -- 275
		"00000000" WHEN "0100010100", -- 276
		"00000000" WHEN "0100010101", -- 277
		"00000000" WHEN "0100010110", -- 278
		"00000000" WHEN "0100010111", -- 279
		"00000000" WHEN "0100011000", -- 280
		"00000000" WHEN "0100011001", -- 281
		"00000000" WHEN "0100011010", -- 282
		"00000000" WHEN "0100011011", -- 283
		"00000000" WHEN "0100011100", -- 284
		"00000000" WHEN "0100011101", -- 285
		"00000000" WHEN "0100011110", -- 286
		"00000000" WHEN "0100011111", -- 287
		"00000000" WHEN "0100100000", -- 288
		"00000011" WHEN "0100100001", -- 289
		"00000000" WHEN "0100100010", -- 290
		"00100110" WHEN "0100100011", -- 291
		"00111111" WHEN "0100100100", -- 292
		"00010110" WHEN "0100100101", -- 293
		"00000000" WHEN "0100100110", -- 294
		"00000000" WHEN "0100100111", -- 295
		"00000000" WHEN "0100101000", -- 296
		"00000000" WHEN "0100101001", -- 297
		"00000000" WHEN "0100101010", -- 298
		"00000000" WHEN "0100101011", -- 299
		"00000000" WHEN "0100101100", -- 300
		"00000000" WHEN "0100101101", -- 301
		"00000000" WHEN "0100101110", -- 302
		"00000000" WHEN "0100101111", -- 303
		"00000000" WHEN "0100110000", -- 304
		"00000000" WHEN "0100110001", -- 305
		"00000000" WHEN "0100110010", -- 306
		"00000000" WHEN "0100110011", -- 307
		"00000000" WHEN "0100110100", -- 308
		"00000000" WHEN "0100110101", -- 309
		"00000000" WHEN "0100110110", -- 310
		"00000000" WHEN "0100110111", -- 311
		"00000000" WHEN "0100111000", -- 312
		"00000000" WHEN "0100111001", -- 313
		"00000000" WHEN "0100111010", -- 314
		"00000000" WHEN "0100111011", -- 315
		"00000000" WHEN "0100111100", -- 316
		"00000000" WHEN "0100111101", -- 317
		"00000000" WHEN "0100111110", -- 318
		"00100010" WHEN "0100111111", -- 319
		"00111111" WHEN "0101000000", -- 320
		"00101111" WHEN "0101000001", -- 321
		"00000000" WHEN "0101000010", -- 322
		"00000000" WHEN "0101000011", -- 323
		"00000000" WHEN "0101000100", -- 324
		"00000000" WHEN "0101000101", -- 325
		"00000000" WHEN "0101000110", -- 326
		"00000000" WHEN "0101000111", -- 327
		"00000000" WHEN "0101001000", -- 328
		"00000000" WHEN "0101001001", -- 329
		"00000000" WHEN "0101001010", -- 330
		"00000000" WHEN "0101001011", -- 331
		"00000000" WHEN "0101001100", -- 332
		"00000000" WHEN "0101001101", -- 333
		"00000000" WHEN "0101001110", -- 334
		"00000000" WHEN "0101001111", -- 335
		"00000000" WHEN "0101010000", -- 336
		"00000000" WHEN "0101010001", -- 337
		"00000000" WHEN "0101010010", -- 338
		"00000000" WHEN "0101010011", -- 339
		"00000000" WHEN "0101010100", -- 340
		"00000000" WHEN "0101010101", -- 341
		"00000000" WHEN "0101010110", -- 342
		"00000000" WHEN "0101010111", -- 343
		"00000000" WHEN "0101011000", -- 344
		"00000000" WHEN "0101011001", -- 345
		"00000000" WHEN "0101011010", -- 346
		"00000010" WHEN "0101011011", -- 347
		"00101111" WHEN "0101011100", -- 348
		"00111111" WHEN "0101011101", -- 349
		"00010001" WHEN "0101011110", -- 350
		"00000000" WHEN "0101011111", -- 351
		"00000000" WHEN "0101100000", -- 352
		"00000000" WHEN "0101100001", -- 353
		"00000000" WHEN "0101100010", -- 354
		"00000000" WHEN "0101100011", -- 355
		"00000000" WHEN "0101100100", -- 356
		"00000000" WHEN "0101100101", -- 357
		"00000000" WHEN "0101100110", -- 358
		"00000000" WHEN "0101100111", -- 359
		"00000000" WHEN "0101101000", -- 360
		"00000000" WHEN "0101101001", -- 361
		"00000000" WHEN "0101101010", -- 362
		"00000000" WHEN "0101101011", -- 363
		"00000000" WHEN "0101101100", -- 364
		"00000000" WHEN "0101101101", -- 365
		"00000000" WHEN "0101101110", -- 366
		"00000000" WHEN "0101101111", -- 367
		"00000000" WHEN "0101110000", -- 368
		"00000000" WHEN "0101110001", -- 369
		"00000000" WHEN "0101110010", -- 370
		"00000000" WHEN "0101110011", -- 371
		"00000000" WHEN "0101110100", -- 372
		"00000000" WHEN "0101110101", -- 373
		"00000000" WHEN "0101110110", -- 374
		"00000000" WHEN "0101110111", -- 375
		"00001000" WHEN "0101111000", -- 376
		"00111100" WHEN "0101111001", -- 377
		"00111000" WHEN "0101111010", -- 378
		"00101000" WHEN "0101111011", -- 379
		"00011011" WHEN "0101111100", -- 380
		"00000000" WHEN "0101111101", -- 381
		"00000000" WHEN "0101111110", -- 382
		"00000000" WHEN "0101111111", -- 383
		"00000000" WHEN "0110000000", -- 384
		"00000000" WHEN "0110000001", -- 385
		"00000000" WHEN "0110000010", -- 386
		"00000000" WHEN "0110000011", -- 387
		"00000000" WHEN "0110000100", -- 388
		"00000000" WHEN "0110000101", -- 389
		"00000000" WHEN "0110000110", -- 390
		"00000000" WHEN "0110000111", -- 391
		"00000000" WHEN "0110001000", -- 392
		"00000000" WHEN "0110001001", -- 393
		"00000000" WHEN "0110001010", -- 394
		"00000000" WHEN "0110001011", -- 395
		"00000000" WHEN "0110001100", -- 396
		"00000000" WHEN "0110001101", -- 397
		"00000000" WHEN "0110001110", -- 398
		"00000000" WHEN "0110001111", -- 399
		"00000000" WHEN "0110010000", -- 400
		"00000000" WHEN "0110010001", -- 401
		"00000000" WHEN "0110010010", -- 402
		"00000000" WHEN "0110010011", -- 403
		"00000000" WHEN "0110010100", -- 404
		"00010100" WHEN "0110010101", -- 405
		"00111100" WHEN "0110010110", -- 406
		"00111111" WHEN "0110010111", -- 407
		"00111111" WHEN "0110011000", -- 408
		"00011101" WHEN "0110011001", -- 409
		"00000110" WHEN "0110011010", -- 410
		"00000000" WHEN "0110011011", -- 411
		"00000000" WHEN "0110011100", -- 412
		"00000000" WHEN "0110011101", -- 413
		"00000000" WHEN "0110011110", -- 414
		"00000000" WHEN "0110011111", -- 415
		"00000000" WHEN "0110100000", -- 416
		"00000000" WHEN "0110100001", -- 417
		"00000000" WHEN "0110100010", -- 418
		"00000000" WHEN "0110100011", -- 419
		"00000000" WHEN "0110100100", -- 420
		"00000000" WHEN "0110100101", -- 421
		"00000000" WHEN "0110100110", -- 422
		"00000000" WHEN "0110100111", -- 423
		"00000000" WHEN "0110101000", -- 424
		"00000000" WHEN "0110101001", -- 425
		"00000000" WHEN "0110101010", -- 426
		"00000000" WHEN "0110101011", -- 427
		"00000000" WHEN "0110101100", -- 428
		"00000000" WHEN "0110101101", -- 429
		"00000000" WHEN "0110101110", -- 430
		"00000000" WHEN "0110101111", -- 431
		"00000000" WHEN "0110110000", -- 432
		"00000000" WHEN "0110110001", -- 433
		"00001011" WHEN "0110110010", -- 434
		"00101110" WHEN "0110110011", -- 435
		"00111111" WHEN "0110110100", -- 436
		"00111111" WHEN "0110110101", -- 437
		"00100101" WHEN "0110110110", -- 438
		"00000110" WHEN "0110110111", -- 439
		"00000000" WHEN "0110111000", -- 440
		"00000000" WHEN "0110111001", -- 441
		"00000000" WHEN "0110111010", -- 442
		"00000000" WHEN "0110111011", -- 443
		"00000000" WHEN "0110111100", -- 444
		"00000000" WHEN "0110111101", -- 445
		"00000000" WHEN "0110111110", -- 446
		"00000000" WHEN "0110111111", -- 447
		"00000000" WHEN "0111000000", -- 448
		"00000000" WHEN "0111000001", -- 449
		"00000000" WHEN "0111000010", -- 450
		"00000000" WHEN "0111000011", -- 451
		"00000000" WHEN "0111000100", -- 452
		"00000000" WHEN "0111000101", -- 453
		"00000000" WHEN "0111000110", -- 454
		"00000000" WHEN "0111000111", -- 455
		"00000000" WHEN "0111001000", -- 456
		"00000000" WHEN "0111001001", -- 457
		"00000000" WHEN "0111001010", -- 458
		"00000000" WHEN "0111001011", -- 459
		"00000000" WHEN "0111001100", -- 460
		"00000000" WHEN "0111001101", -- 461
		"00000000" WHEN "0111001110", -- 462
		"00000100" WHEN "0111001111", -- 463
		"00010111" WHEN "0111010000", -- 464
		"00111111" WHEN "0111010001", -- 465
		"00111111" WHEN "0111010010", -- 466
		"00101110" WHEN "0111010011", -- 467
		"00000000" WHEN "0111010100", -- 468
		"00000000" WHEN "0111010101", -- 469
		"00000000" WHEN "0111010110", -- 470
		"00000000" WHEN "0111010111", -- 471
		"00000000" WHEN "0111011000", -- 472
		"00000000" WHEN "0111011001", -- 473
		"00000000" WHEN "0111011010", -- 474
		"00000000" WHEN "0111011011", -- 475
		"00000000" WHEN "0111011100", -- 476
		"00000000" WHEN "0111011101", -- 477
		"00000000" WHEN "0111011110", -- 478
		"00000000" WHEN "0111011111", -- 479
		"00000000" WHEN "0111100000", -- 480
		"00000000" WHEN "0111100001", -- 481
		"00000000" WHEN "0111100010", -- 482
		"00000000" WHEN "0111100011", -- 483
		"00000000" WHEN "0111100100", -- 484
		"00000000" WHEN "0111100101", -- 485
		"00000000" WHEN "0111100110", -- 486
		"00000000" WHEN "0111100111", -- 487
		"00000000" WHEN "0111101000", -- 488
		"00000000" WHEN "0111101001", -- 489
		"00000000" WHEN "0111101010", -- 490
		"00000000" WHEN "0111101011", -- 491
		"00000000" WHEN "0111101100", -- 492
		"00111110" WHEN "0111101101", -- 493
		"00111111" WHEN "0111101110", -- 494
		"00111110" WHEN "0111101111", -- 495
		"00010000" WHEN "0111110000", -- 496
		"00000000" WHEN "0111110001", -- 497
		"00000000" WHEN "0111110010", -- 498
		"00000000" WHEN "0111110011", -- 499
		"00000000" WHEN "0111110100", -- 500
		"00000000" WHEN "0111110101", -- 501
		"00000000" WHEN "0111110110", -- 502
		"00000000" WHEN "0111110111", -- 503
		"00000000" WHEN "0111111000", -- 504
		"00000000" WHEN "0111111001", -- 505
		"00000000" WHEN "0111111010", -- 506
		"00000000" WHEN "0111111011", -- 507
		"00000000" WHEN "0111111100", -- 508
		"00000000" WHEN "0111111101", -- 509
		"00000000" WHEN "0111111110", -- 510
		"00000000" WHEN "0111111111", -- 511
		"00000000" WHEN "1000000000", -- 512
		"00000000" WHEN "1000000001", -- 513
		"00000000" WHEN "1000000010", -- 514
		"00000000" WHEN "1000000011", -- 515
		"00000000" WHEN "1000000100", -- 516
		"00000000" WHEN "1000000101", -- 517
		"00001011" WHEN "1000000110", -- 518
		"00100000" WHEN "1000000111", -- 519
		"00101101" WHEN "1000001000", -- 520
		"00111111" WHEN "1000001001", -- 521
		"00111111" WHEN "1000001010", -- 522
		"00110011" WHEN "1000001011", -- 523
		"00000000" WHEN "1000001100", -- 524
		"00000000" WHEN "1000001101", -- 525
		"00000000" WHEN "1000001110", -- 526
		"00000000" WHEN "1000001111", -- 527
		"00000000" WHEN "1000010000", -- 528
		"00000000" WHEN "1000010001", -- 529
		"00000000" WHEN "1000010010", -- 530
		"00000000" WHEN "1000010011", -- 531
		"00000000" WHEN "1000010100", -- 532
		"00000000" WHEN "1000010101", -- 533
		"00000000" WHEN "1000010110", -- 534
		"00000000" WHEN "1000010111", -- 535
		"00000000" WHEN "1000011000", -- 536
		"00000000" WHEN "1000011001", -- 537
		"00000000" WHEN "1000011010", -- 538
		"00000000" WHEN "1000011011", -- 539
		"00000000" WHEN "1000011100", -- 540
		"00000000" WHEN "1000011101", -- 541
		"00000000" WHEN "1000011110", -- 542
		"00000000" WHEN "1000011111", -- 543
		"00001001" WHEN "1000100000", -- 544
		"00100101" WHEN "1000100001", -- 545
		"00111001" WHEN "1000100010", -- 546
		"00111111" WHEN "1000100011", -- 547
		"00111111" WHEN "1000100100", -- 548
		"00111111" WHEN "1000100101", -- 549
		"00111110" WHEN "1000100110", -- 550
		"00101101" WHEN "1000100111", -- 551
		"00000000" WHEN "1000101000", -- 552
		"00000000" WHEN "1000101001", -- 553
		"00000000" WHEN "1000101010", -- 554
		"00000000" WHEN "1000101011", -- 555
		"00000000" WHEN "1000101100", -- 556
		"00000000" WHEN "1000101101", -- 557
		"00000000" WHEN "1000101110", -- 558
		"00000000" WHEN "1000101111", -- 559
		"00000000" WHEN "1000110000", -- 560
		"00000000" WHEN "1000110001", -- 561
		"00000000" WHEN "1000110010", -- 562
		"00000000" WHEN "1000110011", -- 563
		"00000000" WHEN "1000110100", -- 564
		"00000000" WHEN "1000110101", -- 565
		"00000000" WHEN "1000110110", -- 566
		"00000000" WHEN "1000110111", -- 567
		"00000000" WHEN "1000111000", -- 568
		"00000000" WHEN "1000111001", -- 569
		"00000110" WHEN "1000111010", -- 570
		"00011100" WHEN "1000111011", -- 571
		"00110111" WHEN "1000111100", -- 572
		"00111111" WHEN "1000111101", -- 573
		"00111111" WHEN "1000111110", -- 574
		"00111111" WHEN "1000111111", -- 575
		"00111111" WHEN "1001000000", -- 576
		"00110010" WHEN "1001000001", -- 577
		"00010011" WHEN "1001000010", -- 578
		"00000000" WHEN "1001000011", -- 579
		"00000000" WHEN "1001000100", -- 580
		"00000000" WHEN "1001000101", -- 581
		"00000000" WHEN "1001000110", -- 582
		"00000000" WHEN "1001000111", -- 583
		"00000000" WHEN "1001001000", -- 584
		"00000000" WHEN "1001001001", -- 585
		"00000000" WHEN "1001001010", -- 586
		"00000000" WHEN "1001001011", -- 587
		"00000000" WHEN "1001001100", -- 588
		"00000000" WHEN "1001001101", -- 589
		"00000000" WHEN "1001001110", -- 590
		"00000000" WHEN "1001001111", -- 591
		"00000000" WHEN "1001010000", -- 592
		"00000000" WHEN "1001010001", -- 593
		"00000000" WHEN "1001010010", -- 594
		"00000000" WHEN "1001010011", -- 595
		"00000101" WHEN "1001010100", -- 596
		"00010000" WHEN "1001010101", -- 597
		"00110101" WHEN "1001010110", -- 598
		"00111111" WHEN "1001010111", -- 599
		"00111111" WHEN "1001011000", -- 600
		"00111111" WHEN "1001011001", -- 601
		"00111111" WHEN "1001011010", -- 602
		"00110001" WHEN "1001011011", -- 603
		"00010100" WHEN "1001011100", -- 604
		"00000000" WHEN "1001011101", -- 605
		"00000000" WHEN "1001011110", -- 606
		"00000000" WHEN "1001011111", -- 607
		"00000000" WHEN "1001100000", -- 608
		"00000000" WHEN "1001100001", -- 609
		"00000000" WHEN "1001100010", -- 610
		"00000000" WHEN "1001100011", -- 611
		"00000000" WHEN "1001100100", -- 612
		"00000000" WHEN "1001100101", -- 613
		"00000000" WHEN "1001100110", -- 614
		"00000000" WHEN "1001100111", -- 615
		"00000000" WHEN "1001101000", -- 616
		"00000000" WHEN "1001101001", -- 617
		"00000000" WHEN "1001101010", -- 618
		"00000000" WHEN "1001101011", -- 619
		"00000000" WHEN "1001101100", -- 620
		"00000000" WHEN "1001101101", -- 621
		"00000100" WHEN "1001101110", -- 622
		"00101010" WHEN "1001101111", -- 623
		"00110110" WHEN "1001110000", -- 624
		"00111111" WHEN "1001110001", -- 625
		"00111111" WHEN "1001110010", -- 626
		"00111111" WHEN "1001110011", -- 627
		"00111111" WHEN "1001110100", -- 628
		"00110000" WHEN "1001110101", -- 629
		"00010100" WHEN "1001110110", -- 630
		"00000010" WHEN "1001110111", -- 631
		"00000000" WHEN "1001111000", -- 632
		"00000000" WHEN "1001111001", -- 633
		"00000000" WHEN "1001111010", -- 634
		"00000000" WHEN "1001111011", -- 635
		"00000000" WHEN "1001111100", -- 636
		"00000000" WHEN "1001111101", -- 637
		"00000000" WHEN "1001111110", -- 638
		"00000000" WHEN "1001111111", -- 639
		"00000000" WHEN "1010000000", -- 640
		"00000000" WHEN "1010000001", -- 641
		"00000000" WHEN "1010000010", -- 642
		"00000000" WHEN "1010000011", -- 643
		"00000000" WHEN "1010000100", -- 644
		"00000000" WHEN "1010000101", -- 645
		"00000000" WHEN "1010000110", -- 646
		"00000000" WHEN "1010000111", -- 647
		"00001101" WHEN "1010001000", -- 648
		"00101011" WHEN "1010001001", -- 649
		"00111000" WHEN "1010001010", -- 650
		"00111111" WHEN "1010001011", -- 651
		"00111111" WHEN "1010001100", -- 652
		"00111111" WHEN "1010001101", -- 653
		"00111111" WHEN "1010001110", -- 654
		"00111101" WHEN "1010001111", -- 655
		"00100001" WHEN "1010010000", -- 656
		"00000010" WHEN "1010010001", -- 657
		"00000000" WHEN "1010010010", -- 658
		"00000000" WHEN "1010010011", -- 659
		"00000000" WHEN "1010010100", -- 660
		"00000000" WHEN "1010010101", -- 661
		"00000000" WHEN "1010010110", -- 662
		"00000000" WHEN "1010010111", -- 663
		"00000000" WHEN "1010011000", -- 664
		"00000000" WHEN "1010011001", -- 665
		"00000000" WHEN "1010011010", -- 666
		"00000000" WHEN "1010011011", -- 667
		"00000000" WHEN "1010011100", -- 668
		"00000000" WHEN "1010011101", -- 669
		"00000000" WHEN "1010011110", -- 670
		"00000000" WHEN "1010011111", -- 671
		"00000000" WHEN "1010100000", -- 672
		"00000000" WHEN "1010100001", -- 673
		"00000000" WHEN "1010100010", -- 674
		"00000000" WHEN "1010100011", -- 675
		"00100010" WHEN "1010100100", -- 676
		"00111111" WHEN "1010100101", -- 677
		"00111111" WHEN "1010100110", -- 678
		"00111111" WHEN "1010100111", -- 679
		"00110101" WHEN "1010101000", -- 680
		"00100001" WHEN "1010101001", -- 681
		"00100001" WHEN "1010101010", -- 682
		"00000100" WHEN "1010101011", -- 683
		"00000000" WHEN "1010101100", -- 684
		"00000000" WHEN "1010101101", -- 685
		"00000000" WHEN "1010101110", -- 686
		"00000000" WHEN "1010101111", -- 687
		"00000000" WHEN "1010110000", -- 688
		"00000000" WHEN "1010110001", -- 689
		"00000000" WHEN "1010110010", -- 690
		"00000000" WHEN "1010110011", -- 691
		"00000000" WHEN "1010110100", -- 692
		"00000000" WHEN "1010110101", -- 693
		"00000000" WHEN "1010110110", -- 694
		"00000000" WHEN "1010110111", -- 695
		"00000000" WHEN "1010111000", -- 696
		"00000000" WHEN "1010111001", -- 697
		"00000000" WHEN "1010111010", -- 698
		"00000000" WHEN "1010111011", -- 699
		"00000000" WHEN "1010111100", -- 700
		"00000000" WHEN "1010111101", -- 701
		"00000000" WHEN "1010111110", -- 702
		"00000000" WHEN "1010111111", -- 703
		"00000000" WHEN "1011000000", -- 704
		"00000000" WHEN "1011000001", -- 705
		"00000000" WHEN "1011000010", -- 706
		"00000000" WHEN "1011000011", -- 707
		"00000000" WHEN "1011000100", -- 708
		"00000000" WHEN "1011000101", -- 709
		"00000000" WHEN "1011000110", -- 710
		"00000000" WHEN "1011000111", -- 711
		"00000000" WHEN "1011001000", -- 712
		"00000000" WHEN "1011001001", -- 713
		"00000000" WHEN "1011001010", -- 714
		"00000000" WHEN "1011001011", -- 715
		"00000000" WHEN "1011001100", -- 716
		"00000000" WHEN "1011001101", -- 717
		"00000000" WHEN "1011001110", -- 718
		"00000000" WHEN "1011001111", -- 719
		"00000000" WHEN "1011010000", -- 720
		"00000000" WHEN "1011010001", -- 721
		"00000000" WHEN "1011010010", -- 722
		"00000000" WHEN "1011010011", -- 723
		"00000000" WHEN "1011010100", -- 724
		"00000000" WHEN "1011010101", -- 725
		"00000000" WHEN "1011010110", -- 726
		"00000000" WHEN "1011010111", -- 727
		"00000000" WHEN "1011011000", -- 728
		"00000000" WHEN "1011011001", -- 729
		"00000000" WHEN "1011011010", -- 730
		"00000000" WHEN "1011011011", -- 731
		"00000000" WHEN "1011011100", -- 732
		"00000000" WHEN "1011011101", -- 733
		"00000000" WHEN "1011011110", -- 734
		"00000000" WHEN "1011011111", -- 735
		"00000000" WHEN "1011100000", -- 736
		"00000000" WHEN "1011100001", -- 737
		"00000000" WHEN "1011100010", -- 738
		"00000000" WHEN "1011100011", -- 739
		"00000000" WHEN "1011100100", -- 740
		"00000000" WHEN "1011100101", -- 741
		"00000000" WHEN "1011100110", -- 742
		"00000000" WHEN "1011100111", -- 743
		"00000000" WHEN "1011101000", -- 744
		"00000000" WHEN "1011101001", -- 745
		"00000000" WHEN "1011101010", -- 746
		"00000000" WHEN "1011101011", -- 747
		"00000000" WHEN "1011101100", -- 748
		"00000000" WHEN "1011101101", -- 749
		"00000000" WHEN "1011101110", -- 750
		"00000000" WHEN "1011101111", -- 751
		"00000000" WHEN "1011110000", -- 752
		"00000000" WHEN "1011110001", -- 753
		"00000000" WHEN "1011110010", -- 754
		"00000000" WHEN "1011110011", -- 755
		"00000000" WHEN "1011110100", -- 756
		"00000000" WHEN "1011110101", -- 757
		"00000000" WHEN "1011110110", -- 758
		"00000000" WHEN "1011110111", -- 759
		"00000000" WHEN "1011111000", -- 760
		"00000000" WHEN "1011111001", -- 761
		"00000000" WHEN "1011111010", -- 762
		"00000000" WHEN "1011111011", -- 763
		"00000000" WHEN "1011111100", -- 764
		"00000000" WHEN "1011111101", -- 765
		"00000000" WHEN "1011111110", -- 766
		"00000000" WHEN "1011111111", -- 767
		"00000000" WHEN "1100000000", -- 768
		"00000000" WHEN "1100000001", -- 769
		"00000000" WHEN "1100000010", -- 770
		"00000000" WHEN "1100000011", -- 771
		"00000000" WHEN "1100000100", -- 772
		"00000000" WHEN "1100000101", -- 773
		"00000000" WHEN "1100000110", -- 774
		"00000000" WHEN "1100000111", -- 775
		"00000000" WHEN "1100001000", -- 776
		"00000000" WHEN "1100001001", -- 777
		"00000000" WHEN "1100001010", -- 778
		"00000000" WHEN "1100001011", -- 779
		"00000000" WHEN "1100001100", -- 780
		"00000000" WHEN "1100001101", -- 781
		"00000000" WHEN "1100001110", -- 782
		"00000000" WHEN "1100001111", -- 783
		"00000000" WHEN OTHERS;
	data_out <= data_out_reg;
END Behavioral;