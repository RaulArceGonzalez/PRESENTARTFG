--------------------------INV------------------------------------
-- This module performs the inverse of the input data (which is the sum of the exponential to perform the softmax function)
---INPUTS
-- data_in : Sum of the exponentials
---OUTPUTS
-- data_out : Inverse of the sum

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE work.tfg_irene_package.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.MATH_REAL.ALL;

ENTITY inverse IS
	PORT (
		data_in : IN STD_LOGIC_VECTOR (input_size_L4fc - 1 DOWNTO 0);
		data_out : OUT STD_LOGIC_VECTOR (input_size_L4fc - 1 DOWNTO 0));
END inverse;

ARCHITECTURE Behavioral OF inverse IS

BEGIN
	WITH data_in SELECT data_out <=
		"11111100" WHEN "10000000",
		"11111011" WHEN "10000001",
		"11111011" WHEN "10000010",
		"11111011" WHEN "10000011",
		"11111011" WHEN "10000100",
		"11111011" WHEN "10000101",
		"11111011" WHEN "10000110",
		"11111011" WHEN "10000111",
		"11111011" WHEN "10001000",
		"11111011" WHEN "10001001",
		"11111011" WHEN "10001010",
		"11111011" WHEN "10001011",
		"11111011" WHEN "10001100",
		"11111011" WHEN "10001101",
		"11111011" WHEN "10001110",
		"11111011" WHEN "10001111",
		"11111011" WHEN "10010000",
		"11111011" WHEN "10010001",
		"11111011" WHEN "10010010",
		"11111011" WHEN "10010011",
		"11111011" WHEN "10010100",
		"11111011" WHEN "10010101",
		"11111011" WHEN "10010110",
		"11111011" WHEN "10010111",
		"11111011" WHEN "10011000",
		"11111011" WHEN "10011001",
		"11111010" WHEN "10011010",
		"11111010" WHEN "10011011",
		"11111010" WHEN "10011100",
		"11111010" WHEN "10011101",
		"11111010" WHEN "10011110",
		"11111010" WHEN "10011111",
		"11111010" WHEN "10100000",
		"11111010" WHEN "10100001",
		"11111010" WHEN "10100010",
		"11111010" WHEN "10100011",
		"11111010" WHEN "10100100",
		"11111010" WHEN "10100101",
		"11111010" WHEN "10100110",
		"11111010" WHEN "10100111",
		"11111010" WHEN "10101000",
		"11111010" WHEN "10101001",
		"11111010" WHEN "10101010",
		"11111001" WHEN "10101011",
		"11111001" WHEN "10101100",
		"11111001" WHEN "10101101",
		"11111001" WHEN "10101110",
		"11111001" WHEN "10101111",
		"11111001" WHEN "10110000",
		"11111001" WHEN "10110001",
		"11111001" WHEN "10110010",
		"11111001" WHEN "10110011",
		"11111001" WHEN "10110100",
		"11111001" WHEN "10110101",
		"11111001" WHEN "10110110",
		"11111000" WHEN "10110111",
		"11111000" WHEN "10111000",
		"11111000" WHEN "10111001",
		"11111000" WHEN "10111010",
		"11111000" WHEN "10111011",
		"11111000" WHEN "10111100",
		"11111000" WHEN "10111101",
		"11111000" WHEN "10111110",
		"11111000" WHEN "10111111",
		"11111000" WHEN "11000000",
		"11110111" WHEN "11000001",
		"11110111" WHEN "11000010",
		"11110111" WHEN "11000011",
		"11110111" WHEN "11000100",
		"11110111" WHEN "11000101",
		"11110111" WHEN "11000110",
		"11110111" WHEN "11000111",
		"11110110" WHEN "11001000",
		"11110110" WHEN "11001001",
		"11110110" WHEN "11001010",
		"11110110" WHEN "11001011",
		"11110110" WHEN "11001100",
		"11110101" WHEN "11001101",
		"11110101" WHEN "11001110",
		"11110101" WHEN "11001111",
		"11110101" WHEN "11010000",
		"11110101" WHEN "11010001",
		"11110100" WHEN "11010010",
		"11110100" WHEN "11010011",
		"11110100" WHEN "11010100",
		"11110100" WHEN "11010101",
		"11110011" WHEN "11010110",
		"11110011" WHEN "11010111",
		"11110011" WHEN "11011000",
		"11110010" WHEN "11011001",
		"11110010" WHEN "11011010",
		"11110010" WHEN "11011011",
		"11110001" WHEN "11011100",
		"11110001" WHEN "11011101",
		"11110000" WHEN "11011110",
		"11110000" WHEN "11011111",
		"11110000" WHEN "11100000",
		"11101111" WHEN "11100001",
		"11101110" WHEN "11100010",
		"11101110" WHEN "11100011",
		"11101101" WHEN "11100100",
		"11101101" WHEN "11100101",
		"11101100" WHEN "11100110",
		"11101011" WHEN "11100111",
		"11101010" WHEN "11101000",
		"11101001" WHEN "11101001",
		"11101000" WHEN "11101010",
		"11100111" WHEN "11101011",
		"11100110" WHEN "11101100",
		"11100101" WHEN "11101101",
		"11100011" WHEN "11101110",
		"11100001" WHEN "11101111",
		"11100000" WHEN "11110000",
		"11011101" WHEN "11110001",
		"11011011" WHEN "11110010",
		"11011000" WHEN "11110011",
		"11010101" WHEN "11110100",
		"11010001" WHEN "11110101",
		"11001100" WHEN "11110110",
		"11000111" WHEN "11110111",
		"11000000" WHEN "11111000",
		"10110110" WHEN "11111001",
		"10101010" WHEN "11111010",
		"10011001" WHEN "11111011",
		"10000000" WHEN "11111100",
		"10000000" WHEN "11111101",
		"10000000" WHEN "11111110",
		"10000000" WHEN "11111111",
		"01111111" WHEN "00000000",
		"01111111" WHEN "00000001",
		"01111111" WHEN "00000010",
		"01111111" WHEN "00000011",
		"01111111" WHEN "00000100",
		"01100110" WHEN "00000101",
		"01010101" WHEN "00000110",
		"01001001" WHEN "00000111",
		"01000000" WHEN "00001000",
		"00111000" WHEN "00001001",
		"00110011" WHEN "00001010",
		"00101110" WHEN "00001011",
		"00101010" WHEN "00001100",
		"00100111" WHEN "00001101",
		"00100100" WHEN "00001110",
		"00100010" WHEN "00001111",
		"00100000" WHEN "00010000",
		"00011110" WHEN "00010001",
		"00011100" WHEN "00010010",
		"00011010" WHEN "00010011",
		"00011001" WHEN "00010100",
		"00011000" WHEN "00010101",
		"00010111" WHEN "00010110",
		"00010110" WHEN "00010111",
		"00010101" WHEN "00011000",
		"00010100" WHEN "00011001",
		"00010011" WHEN "00011010",
		"00010010" WHEN "00011011",
		"00010010" WHEN "00011100",
		"00010001" WHEN "00011101",
		"00010001" WHEN "00011110",
		"00010000" WHEN "00011111",
		"00010000" WHEN "00100000",
		"00001111" WHEN "00100001",
		"00001111" WHEN "00100010",
		"00001110" WHEN "00100011",
		"00001110" WHEN "00100100",
		"00001101" WHEN "00100101",
		"00001101" WHEN "00100110",
		"00001101" WHEN "00100111",
		"00001100" WHEN "00101000",
		"00001100" WHEN "00101001",
		"00001100" WHEN "00101010",
		"00001011" WHEN "00101011",
		"00001011" WHEN "00101100",
		"00001011" WHEN "00101101",
		"00001011" WHEN "00101110",
		"00001010" WHEN "00101111",
		"00001010" WHEN "00110000",
		"00001010" WHEN "00110001",
		"00001010" WHEN "00110010",
		"00001010" WHEN "00110011",
		"00001001" WHEN "00110100",
		"00001001" WHEN "00110101",
		"00001001" WHEN "00110110",
		"00001001" WHEN "00110111",
		"00001001" WHEN "00111000",
		"00001000" WHEN "00111001",
		"00001000" WHEN "00111010",
		"00001000" WHEN "00111011",
		"00001000" WHEN "00111100",
		"00001000" WHEN "00111101",
		"00001000" WHEN "00111110",
		"00001000" WHEN "00111111",
		"00001000" WHEN "01000000",
		"00000111" WHEN "01000001",
		"00000111" WHEN "01000010",
		"00000111" WHEN "01000011",
		"00000111" WHEN "01000100",
		"00000111" WHEN "01000101",
		"00000111" WHEN "01000110",
		"00000111" WHEN "01000111",
		"00000111" WHEN "01001000",
		"00000111" WHEN "01001001",
		"00000110" WHEN "01001010",
		"00000110" WHEN "01001011",
		"00000110" WHEN "01001100",
		"00000110" WHEN "01001101",
		"00000110" WHEN "01001110",
		"00000110" WHEN "01001111",
		"00000110" WHEN "01010000",
		"00000110" WHEN "01010001",
		"00000110" WHEN "01010010",
		"00000110" WHEN "01010011",
		"00000110" WHEN "01010100",
		"00000110" WHEN "01010101",
		"00000101" WHEN "01010110",
		"00000101" WHEN "01010111",
		"00000101" WHEN "01011000",
		"00000101" WHEN "01011001",
		"00000101" WHEN "01011010",
		"00000101" WHEN "01011011",
		"00000101" WHEN "01011100",
		"00000101" WHEN "01011101",
		"00000101" WHEN "01011110",
		"00000101" WHEN "01011111",
		"00000101" WHEN "01100000",
		"00000101" WHEN "01100001",
		"00000101" WHEN "01100010",
		"00000101" WHEN "01100011",
		"00000101" WHEN "01100100",
		"00000101" WHEN "01100101",
		"00000101" WHEN "01100110",
		"00000100" WHEN "01100111",
		"00000100" WHEN "01101000",
		"00000100" WHEN "01101001",
		"00000100" WHEN "01101010",
		"00000100" WHEN "01101011",
		"00000100" WHEN "01101100",
		"00000100" WHEN "01101101",
		"00000100" WHEN "01101110",
		"00000100" WHEN "01101111",
		"00000100" WHEN "01110000",
		"00000100" WHEN "01110001",
		"00000100" WHEN "01110010",
		"00000100" WHEN "01110011",
		"00000100" WHEN "01110100",
		"00000100" WHEN "01110101",
		"00000100" WHEN "01110110",
		"00000100" WHEN "01110111",
		"00000100" WHEN "01111000",
		"00000100" WHEN "01111001",
		"00000100" WHEN "01111010",
		"00000100" WHEN "01111011",
		"00000100" WHEN "01111100",
		"00000100" WHEN "01111101",
		"00000100" WHEN "01111110",
		"00000100" WHEN "01111111",
		"00000000" WHEN OTHERS;
END Behavioral;