--------------------------Sigmoid------------------------------------
-- This module performs the sigmoid function with a LUT
---INPUTS
-- data_in : Results of the convolution operations.
---OUTPUTS
-- data_out : Sigmoid of the input data.

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE work.tfg_irene_package.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.MATH_REAL.ALL;

ENTITY sigmoid_L3 IS
	PORT (
		data_in : IN STD_LOGIC_VECTOR(input_sizeL3 - 1 DOWNTO 0);
		data_out : OUT STD_LOGIC_VECTOR(input_sizeL3 - 1 DOWNTO 0));
END sigmoid_L3;

ARCHITECTURE Behavioral OF sigmoid_L3 IS

BEGIN
	WITH data_in SELECT data_out <=
		"00000111" WHEN "10000000",
		"00000111" WHEN "10000001",
		"00000111" WHEN "10000010",
		"00000111" WHEN "10000011",
		"00001000" WHEN "10000100",
		"00001000" WHEN "10000101",
		"00001000" WHEN "10000110",
		"00001000" WHEN "10000111",
		"00001000" WHEN "10001000",
		"00001000" WHEN "10001001",
		"00001000" WHEN "10001010",
		"00001000" WHEN "10001011",
		"00001000" WHEN "10001100",
		"00001001" WHEN "10001101",
		"00001001" WHEN "10001110",
		"00001001" WHEN "10001111",
		"00001001" WHEN "10010000",
		"00001001" WHEN "10010001",
		"00001001" WHEN "10010010",
		"00001001" WHEN "10010011",
		"00001001" WHEN "10010100",
		"00001010" WHEN "10010101",
		"00001010" WHEN "10010110",
		"00001010" WHEN "10010111",
		"00001010" WHEN "10011000",
		"00001010" WHEN "10011001",
		"00001010" WHEN "10011010",
		"00001010" WHEN "10011011",
		"00001011" WHEN "10011100",
		"00001011" WHEN "10011101",
		"00001011" WHEN "10011110",
		"00001011" WHEN "10011111",
		"00001011" WHEN "10100000",
		"00001011" WHEN "10100001",
		"00001011" WHEN "10100010",
		"00001100" WHEN "10100011",
		"00001100" WHEN "10100100",
		"00001100" WHEN "10100101",
		"00001100" WHEN "10100110",
		"00001100" WHEN "10100111",
		"00001100" WHEN "10101000",
		"00001101" WHEN "10101001",
		"00001101" WHEN "10101010",
		"00001101" WHEN "10101011",
		"00001101" WHEN "10101100",
		"00001101" WHEN "10101101",
		"00001101" WHEN "10101110",
		"00001110" WHEN "10101111",
		"00001110" WHEN "10110000",
		"00001110" WHEN "10110001",
		"00001110" WHEN "10110010",
		"00001110" WHEN "10110011",
		"00001110" WHEN "10110100",
		"00001111" WHEN "10110101",
		"00001111" WHEN "10110110",
		"00001111" WHEN "10110111",
		"00001111" WHEN "10111000",
		"00001111" WHEN "10111001",
		"00010000" WHEN "10111010",
		"00010000" WHEN "10111011",
		"00010000" WHEN "10111100",
		"00010000" WHEN "10111101",
		"00010000" WHEN "10111110",
		"00010001" WHEN "10111111",
		"00010001" WHEN "11000000",
		"00010001" WHEN "11000001",
		"00010001" WHEN "11000010",
		"00010001" WHEN "11000011",
		"00010010" WHEN "11000100",
		"00010010" WHEN "11000101",
		"00010010" WHEN "11000110",
		"00010010" WHEN "11000111",
		"00010010" WHEN "11001000",
		"00010011" WHEN "11001001",
		"00010011" WHEN "11001010",
		"00010011" WHEN "11001011",
		"00010011" WHEN "11001100",
		"00010011" WHEN "11001101",
		"00010100" WHEN "11001110",
		"00010100" WHEN "11001111",
		"00010100" WHEN "11010000",
		"00010100" WHEN "11010001",
		"00010100" WHEN "11010010",
		"00010101" WHEN "11010011",
		"00010101" WHEN "11010100",
		"00010101" WHEN "11010101",
		"00010101" WHEN "11010110",
		"00010110" WHEN "11010111",
		"00010110" WHEN "11011000",
		"00010110" WHEN "11011001",
		"00010110" WHEN "11011010",
		"00010110" WHEN "11011011",
		"00010111" WHEN "11011100",
		"00010111" WHEN "11011101",
		"00010111" WHEN "11011110",
		"00010111" WHEN "11011111",
		"00011000" WHEN "11100000",
		"00011000" WHEN "11100001",
		"00011000" WHEN "11100010",
		"00011000" WHEN "11100011",
		"00011001" WHEN "11100100",
		"00011001" WHEN "11100101",
		"00011001" WHEN "11100110",
		"00011001" WHEN "11100111",
		"00011010" WHEN "11101000",
		"00011010" WHEN "11101001",
		"00011010" WHEN "11101010",
		"00011010" WHEN "11101011",
		"00011011" WHEN "11101100",
		"00011011" WHEN "11101101",
		"00011011" WHEN "11101110",
		"00011011" WHEN "11101111",
		"00011100" WHEN "11110000",
		"00011100" WHEN "11110001",
		"00011100" WHEN "11110010",
		"00011100" WHEN "11110011",
		"00011101" WHEN "11110100",
		"00011101" WHEN "11110101",
		"00011101" WHEN "11110110",
		"00011101" WHEN "11110111",
		"00011110" WHEN "11111000",
		"00011110" WHEN "11111001",
		"00011110" WHEN "11111010",
		"00011110" WHEN "11111011",
		"00011111" WHEN "11111100",
		"00011111" WHEN "11111101",
		"00011111" WHEN "11111110",
		"00011111" WHEN "11111111",
		"00100000" WHEN "00000000",
		"00100000" WHEN "00000001",
		"00100000" WHEN "00000010",
		"00100000" WHEN "00000011",
		"00100000" WHEN "00000100",
		"00100001" WHEN "00000101",
		"00100001" WHEN "00000110",
		"00100001" WHEN "00000111",
		"00100001" WHEN "00001000",
		"00100010" WHEN "00001001",
		"00100010" WHEN "00001010",
		"00100010" WHEN "00001011",
		"00100010" WHEN "00001100",
		"00100011" WHEN "00001101",
		"00100011" WHEN "00001110",
		"00100011" WHEN "00001111",
		"00100011" WHEN "00010000",
		"00100100" WHEN "00010001",
		"00100100" WHEN "00010010",
		"00100100" WHEN "00010011",
		"00100100" WHEN "00010100",
		"00100101" WHEN "00010101",
		"00100101" WHEN "00010110",
		"00100101" WHEN "00010111",
		"00100101" WHEN "00011000",
		"00100110" WHEN "00011001",
		"00100110" WHEN "00011010",
		"00100110" WHEN "00011011",
		"00100110" WHEN "00011100",
		"00100111" WHEN "00011101",
		"00100111" WHEN "00011110",
		"00100111" WHEN "00011111",
		"00100111" WHEN "00100000",
		"00101000" WHEN "00100001",
		"00101000" WHEN "00100010",
		"00101000" WHEN "00100011",
		"00101000" WHEN "00100100",
		"00101001" WHEN "00100101",
		"00101001" WHEN "00100110",
		"00101001" WHEN "00100111",
		"00101001" WHEN "00101000",
		"00101001" WHEN "00101001",
		"00101010" WHEN "00101010",
		"00101010" WHEN "00101011",
		"00101010" WHEN "00101100",
		"00101010" WHEN "00101101",
		"00101011" WHEN "00101110",
		"00101011" WHEN "00101111",
		"00101011" WHEN "00110000",
		"00101011" WHEN "00110001",
		"00101011" WHEN "00110010",
		"00101100" WHEN "00110011",
		"00101100" WHEN "00110100",
		"00101100" WHEN "00110101",
		"00101100" WHEN "00110110",
		"00101100" WHEN "00110111",
		"00101101" WHEN "00111000",
		"00101101" WHEN "00111001",
		"00101101" WHEN "00111010",
		"00101101" WHEN "00111011",
		"00101101" WHEN "00111100",
		"00101110" WHEN "00111101",
		"00101110" WHEN "00111110",
		"00101110" WHEN "00111111",
		"00101110" WHEN "01000000",
		"00101110" WHEN "01000001",
		"00101111" WHEN "01000010",
		"00101111" WHEN "01000011",
		"00101111" WHEN "01000100",
		"00101111" WHEN "01000101",
		"00101111" WHEN "01000110",
		"00110000" WHEN "01000111",
		"00110000" WHEN "01001000",
		"00110000" WHEN "01001001",
		"00110000" WHEN "01001010",
		"00110000" WHEN "01001011",
		"00110001" WHEN "01001100",
		"00110001" WHEN "01001101",
		"00110001" WHEN "01001110",
		"00110001" WHEN "01001111",
		"00110001" WHEN "01010000",
		"00110001" WHEN "01010001",
		"00110010" WHEN "01010010",
		"00110010" WHEN "01010011",
		"00110010" WHEN "01010100",
		"00110010" WHEN "01010101",
		"00110010" WHEN "01010110",
		"00110010" WHEN "01010111",
		"00110011" WHEN "01011000",
		"00110011" WHEN "01011001",
		"00110011" WHEN "01011010",
		"00110011" WHEN "01011011",
		"00110011" WHEN "01011100",
		"00110011" WHEN "01011101",
		"00110100" WHEN "01011110",
		"00110100" WHEN "01011111",
		"00110100" WHEN "01100000",
		"00110100" WHEN "01100001",
		"00110100" WHEN "01100010",
		"00110100" WHEN "01100011",
		"00110100" WHEN "01100100",
		"00110101" WHEN "01100101",
		"00110101" WHEN "01100110",
		"00110101" WHEN "01100111",
		"00110101" WHEN "01101000",
		"00110101" WHEN "01101001",
		"00110101" WHEN "01101010",
		"00110101" WHEN "01101011",
		"00110110" WHEN "01101100",
		"00110110" WHEN "01101101",
		"00110110" WHEN "01101110",
		"00110110" WHEN "01101111",
		"00110110" WHEN "01110000",
		"00110110" WHEN "01110001",
		"00110110" WHEN "01110010",
		"00110110" WHEN "01110011",
		"00110111" WHEN "01110100",
		"00110111" WHEN "01110101",
		"00110111" WHEN "01110110",
		"00110111" WHEN "01110111",
		"00110111" WHEN "01111000",
		"00110111" WHEN "01111001",
		"00110111" WHEN "01111010",
		"00110111" WHEN "01111011",
		"00110111" WHEN "01111100",
		"00111000" WHEN "01111101",
		"00111000" WHEN "01111110",
		"00111000" WHEN "01111111",
		"00000000" WHEN OTHERS;
END Behavioral;